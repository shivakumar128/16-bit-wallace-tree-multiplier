`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:19:13 02/29/2020 
// Design Name: 
// Module Name:    muull 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:09:34 02/28/2020 
// Design Name: 
// Module Name:    multiplexer 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module multiplier(out1,of,out2,a,b
    );
	 output [15:0]out1,out2;
	 input [15:0]a,b;
	 output of;
	 wire [15:0] p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15;
	 wire s11,s12,s13,s14,s16,s17,s18,s19,s110,s111,s112,s113,s114,s115,s21,s22,s23,s24,s25,s26,s27,s28,s29,s210,s211,s212,s213,s214,s215,
	 s31,s32,s33,s34,s35,s36,s37,s38,s39,s310,s311,s312,s313,s314,s315,s41,s42,s43,s44,s45,s46,s47,s48,s49,s410,s411,s412,s413,s414,s415,
	s15,s52,s53,s54,s55,s56,s57,s58,s59,s510,s511,s512,s513,s514,s515,s61,s62,s63,s64,s65,s66,s67,s68,s69,s610,s611,s612,s613,s614,s615,
	s71,s72,s73,s74,s75,s76,s77,s78,s79,s710,s711,s712,s713,s714,s715,s81,s82,s83,s84,s85,s86,s87,s88,s89,s810,s811,s812,s813,s814,s815,
	s91,s92,s93,s94,s95,s96,s97,s98,s99,s910,s911,s912,s913,s914,s915,s101,s102,s103,s104,s105,s106,s107,s108,s109,s1010,s1011,s1012,s1013,s1014,s1015,
	s11_1,s11_2,s11_3,s11_4,s11_5,s116,s117,s118,s119,s1110,s1111,s1112,s1113,s1114,s1115,s121,s122,s123,s124,s125,s126,s127,s128,s129,s1210,s1211,s1212,s1213,s1214,s1215,
	s131,s132,s133,s134,s135,s136,s137,s138,s139,s1310,s1311,s1312,s1313,s1314,s1315,s141,s142,s143,s144,s145,s146,s147,s148,s149,s1410,s1411,s1412,s1413,s1414,s1415;
	
	
	
	//first stage
	wire c11,cc1,c12,c13,c14,c16,c17,c18,c19,c110,c111,c112,c113,c114,c115,c116,c21,c22,c23,c24,c25,c26,c27,c28,c29,c210,c211,c212,c213,c214,c215,c216,
	 c31,c32,c33,c34,c35,c36,c37,c38,c39,c310,c311,c312,c313,c314,c315,c316,c41,c42,c43,c44,c45,c46,c47,c48,c49,c410,c411,c412,c413,c414,c415,c416,
	c15,c52,c53,c54,c55,c56,c57,c58,c59,c510,c511,c512,c513,c514,c515,c516,c61,c62,c63,c64,c65,c66,c67,c68,c69,c610,c611,c612,c613,c614,c615,c616,
	c71,c72,c73,c74,c75,c76,c77,c78,c79,c710,c711,c712,c713,c714,c715,c716,c81,c82,c83,c84,c85,c86,c87,c88,c89,c810,c811,c812,c813,c814,c815,c816,
	c91,c92,c93,c94,c95,c96,c97,c98,c99,c910,c911,c912,c913,c914,c915,c916,c101,c102,c103,c104,c105,c106,c107,c108,c109,c1010,c1011,c1012,c1013,c1014,c1015,c1016,
	c11_1,c11_2,c11_3,c11_4,c11_5,c11_6,c117,c118,c119,c1110,c1111,c1112,c1113,c1114,c1115,c1116,c121,c122,c123,c124,c125,c126,c127,c128,c129,c1210,c1211,c1212,c1213,c1214,c1215,c1216,
	c131,c132,c133,c134,c135,c136,c137,c138,c139,c1310,c1311,c1312,c1313,c1314,c1315,c1316,c141,c142,c143,c144,c145,c146,c147,c148,c149,c1410,c1411,c1412,c1413,c1414,c1415,c1416,c151,c152,c153,c154,c155,c156,c157,c158,c159,c1510,c1511,c1512,c1513,c1514,c1515,c1516,c1517;
	

	 assign p0=a & {16{b[0]}};
	 assign p1=a & {16{b[1]}};
	 assign p2=a & {16{b[2]}};
	 assign p3=a & {16{b[3]}};
	 assign p4=a & {16{b[4]}};
	 assign p5=a & {16{b[5]}};
	 assign p6=a & {16{b[6]}};
	 assign p7=a & {16{b[7]}};
	 assign p8=a & {16{b[8]}};
	 assign p9=a & {16{b[9]}};
	 assign p10=a & {16{b[10]}};
	 assign p11=a & {16{b[11]}};
	 assign p12=a & {16{b[12]}};
	 assign p13=a & {16{b[13]}};
	 assign p14=a & {16{b[14]}};
	 assign p15=a & {16{b[15]}};
	 assign out1[0]=p0[0];
	ha h1(out1[1],c11,p0[1],p1[0]);
	fa f1(s11,c12,p0[2],p1[1],p2[0]);
	fa f2(s12,c13,p0[3],p1[2],p2[1]);
	fa f3(s13,c14,p0[4],p1[3],p2[2]);
	fa f4(s14,c15,p0[5],p1[4],p2[3]);
	fa f5(s15,c16,p0[6],p1[5],p2[4]);
	fa f6(s16,c17,p0[7],p1[6],p2[5]);
	fa f7(s17,c18,p0[8],p1[7],p2[6]);
	fa f8(s18,c19,p0[9],p1[8],p2[7]);
	fa f9(s19,c110,p0[10],p1[9],p2[8]);
	fa f10(s110,c111,p0[11],p1[10],p2[9]);
	fa f11(s111,c112,p0[12],p1[11],p2[10]);
	fa f12(s112,c113,p0[13],p1[12],p2[11]);
	fa f13(s113,c114,p0[14],p1[13],p2[12]);
	fa f111(s114,c115,p0[15],p1[14],p2[13]);
	ha h2(s115,c116,p1[15],p2[14]);
	//second stage
	ha h3(out1[2],c21,s11,c11);
	fa f14(s21,c22,s12,c12,p3[0]);
	fa f15(s22,c23,s13,c13,p3[1]);
	fa f16(s23,c24,s14,c14,p3[2]);
	fa f17(s24,c25,s15,c15,p3[3]);
	fa f18(s25,c26,s16,c16,p3[4]);
	fa f19(s26,c27,s17,c17,p3[5]);
	fa f20(s27,c28,s18,c18,p3[6]);
	fa f21(s28,c29,s19,c19,p3[7]);
	fa f22(s29,c210,s110,c110,p3[8]);
	fa f23(s210,c211,s111,c111,p3[9]);
	fa f24(s211,c212,s112,c112,p3[10]);
	fa f25(s212,c213,s113,c113,p3[11]);
	fa f26(s213,c214,s114,c114,p3[12]);
	fa f27(s214,c215,s115,c115,p3[13]);
	fa h4(s215,c216,p2[15],p3[14],c116);
	//stage three
	ha h5(out1[3],c31,s21,c21);
	fa f28(s31,c32,s22,c22,p4[0]);
	fa f29(s32,c33,s23,c23,p4[1]);
	fa f30(s33,c34,s24,c24,p4[2]);
	fa f31(s34,c35,s25,c25,p4[3]);
	fa f32(s35,c36,s26,c26,p4[4]);
	fa f33(s36,c37,s27,c27,p4[5]);
	fa f34(s37,c38,s28,c28,p4[6]);
	fa f35(s38,c39,s29,c29,p4[7]);
	fa f36(s39,c310,s210,c210,p4[8]);
	fa f37(s310,c311,s211,c211,p4[9]);
	fa f38(s311,c312,s212,c212,p4[10]);
	fa f39(s312,c313,s213,c213,p4[11]);
	fa f40(s313,c314,s214,c214,p4[12]);
	fa f41(s314,c315,s215,c215,p4[13]);
	fa h6(s315,c316,p3[15],p4[14],c216);
	//stage four
	ha h7(out1[4],c41,s31,c31);
	fa f42(s41,c42,s32,c32,p4[0]);
	fa f43(s42,c43,s33,c33,p4[1]);
	fa f44(s43,c44,s34,c34,p4[2]);
	fa f45(s44,c45,s35,c35,p4[3]);
	fa f46(s45,c46,s36,c36,p4[4]);
	fa f47(s46,c47,s37,c37,p4[5]);
	fa f48(s47,c48,s38,c38,p4[6]);
	fa f49(s48,c49,s39,c39,p4[7]);
	fa f50(s49,c410,s310,c310,p4[8]);
	fa f51(s410,c411,s311,c311,p4[9]);
	fa f52(s411,c412,s312,c312,p4[10]);
	fa f53(s412,c413,s313,c313,p4[11]);
	fa f54(s413,c414,s314,c314,p4[12]);
	fa f55(s414,c415,s315,c315,p4[13]);
	fa h8(s415,c416,p4[15],p5[14],c316);
	//stage five
	ha h9(out1[5],c51,s41,c41);
	fa f56(s51,c52,s42,c42,p5[0]);
	fa f57(s52,c53,s43,c43,p5[1]);
	fa f58(s53,c54,s44,c44,p5[2]);
	fa f59(s54,c55,s45,c45,p5[3]);
	fa f60(s55,c56,s46,c46,p5[4]);
	fa f61(s56,c57,s47,c47,p5[5]);
	fa f62(s57,c58,s48,c48,p5[6]);
	fa f63(s58,c59,s49,c49,p5[7]);
	fa f64(s59,c510,s410,c410,p5[8]);
	fa f65(s510,c511,s411,c411,p5[9]);
	fa f66(s511,c512,s412,c412,p5[10]);
	fa f67(s512,c513,s413,c413,p5[11]);
	fa f68(s513,c514,s414,c414,p5[12]);
	fa f69(s514,c515,s415,c415,p5[13]);
	fa h10(s515,c516,p5[15],p6[14],c416);
	//stage 6
	ha h11(out1[6],c61,s51,c51);
	fa f70(s61,c62,s52,c52,p7[0]);
	fa f71(s62,c63,s53,c53,p7[1]);
	fa f72(s63,c64,s54,c54,p7[2]);
	fa f73(s64,c65,s55,c55,p7[3]);
	fa f74(s65,c66,s56,c56,p7[4]);
	fa f75(s66,c67,s57,c57,p7[5]);
	fa f76(s67,c68,s58,c58,p7[6]);
	fa f77(s68,c69,s59,c59,p7[7]);
	fa f78(s69,c610,s510,c510,p7[8]);
	fa f79(s610,c611,s511,c511,p7[9]);
	fa f80(s611,c612,s512,c512,p7[10]);
	fa f81(s612,c613,s513,c513,p7[11]);
	fa f82(s613,c614,s514,c514,p7[12]);
	fa f83(s614,c615,s515,c515,p7[13]);
	fa h12(s615,c616,p6[15],p7[14],c516);
	//stage 7
	ha h13(out1[7],c71,s61,c61);
	fa f84(s71,c72,s62,c62,p8[0]);
	fa f85(s72,c73,s63,c63,p8[1]);
	fa f86(s73,c74,s64,c64,p8[2]);
	fa f87(s74,c75,s65,c65,p8[3]);
	fa f88(s75,c76,s66,c66,p8[4]);
	fa f89(s76,c77,s67,c67,p8[5]);
	fa f90(s77,c78,s68,c68,p8[6]);
	fa f91(s78,c79,s69,c69,p8[7]);
	fa f92(s79,c710,s610,c610,p8[8]);
	fa f93(s710,c711,s611,c611,p8[9]);
	fa f94(s711,c712,s612,c612,p8[10]);
	fa f95(s712,c713,s613,c613,p8[11]);
	fa f96(s713,c714,s614,c614,p8[12]);
	fa f97(s714,c715,s615,c615,p8[13]);
	fa h14(s715,c716,p7[15],p8[14],c616);
	//stage 8
	ha h15(out1[8],c81,s71,c71);
	fa f98(s81,c82,s72,c72,p9[0]);
	fa f99(s82,c83,s73,c73,p9[1]);
	fa f100(s83,c84,s74,c74,p9[2]);
	fa f101(s84,c85,s75,c75,p9[3]);
	fa f102(s85,c86,s76,c76,p9[4]);
	fa f103(s86,c87,s77,c77,p9[5]);
	fa f104(s87,c88,s78,c78,p9[6]);
	fa f105(s88,c89,s79,c79,p9[7]);
	fa f106(s89,c810,s710,c710,p9[8]);
	fa f107(s810,c811,s711,c711,p9[9]);
	fa f108(s811,c812,s712,c712,p9[10]);
	fa f109(s812,c813,s713,c713,p9[11]);
	fa f110(s813,c814,s714,c714,p9[12]);
	fa f1111(s814,c815,s715,c715,p9[13]);
	fa h16(s815,c816,p8[15],p9[14],c716);
	//stage 9
	ha h17(out1[9],c91,s81,c81);
	fa f112(s91,c92,s82,c82,p10[0]);
	fa f113(s92,c93,s83,c83,p10[1]);
	fa f114(s93,c94,s84,c84,p10[2]);
	fa f115(s94,c95,s85,c85,p10[3]);
	fa f116(s95,c96,s86,c86,p10[4]);
	fa f117(s96,c97,s87,c87,p10[5]);
	fa f118(s97,c98,s88,c88,p10[6]);
	fa f119(s98,c99,s89,c89,p10[7]);
	fa f120(s99,c910,s810,c810,p10[8]);
	fa f121(s910,c911,s811,c811,p10[9]);
	fa f122(s911,c912,s812,c812,p10[10]);
	fa f123(s912,c913,s813,c813,p10[11]);
	fa f124(s913,c914,s814,c814,p10[12]);
	fa f125(s914,c915,s815,c815,p10[13]);
	fa h18(s915,c916,p9[15],p10[14],c816);
	//stage 10
	ha h19(out1[10],c101,s91,c91);
	fa f126(s101,c102,s92,c92,p11[0]);
	fa f127(s102,c103,s93,c93,p11[1]);
	fa f128(s103,c104,s94,c94,p11[2]);
	fa f129(s104,c105,s95,c95,p11[3]);
	fa f130(s105,c106,s96,c96,p11[4]);
	fa f131(s106,c107,s97,c97,p11[5]);
	fa f132(s107,c108,s98,c98,p11[6]);
	fa f133(s108,c109,s99,c99,p11[7]);
	fa f134(s109,c1010,s910,c910,p11[8]);
	fa f135(s1010,c1011,s911,c911,p11[9]);
	fa f136(s1011,c1012,s912,c912,p11[10]);
	fa f137(s1012,c1013,s913,c913,p11[11]);
	fa f138(s1013,c1014,s914,c914,p11[12]);
	fa f139(s1014,c1015,s915,c915,p11[13]);
	fa h20(s1015,c1016,p10[15],p11[14],c916);
	//stage 11
	ha h21(out1[11],c11_1,s101,c101);
	fa f140(s11_1,c11_2,s102,c102,p12[0]);
	fa f141(s11_2,c11_3,s103,c103,p12[1]);
	fa f142(s11_3,c11_4,s104,c104,p12[2]);
	fa f143(s11_4,c11_5,s105,c105,p12[3]);
	fa f144(s11_5,c11_6,s106,c106,p12[4]);
	fa f145(s116,c117,s107,c107,p12[5]);
	fa f146(s117,c118,s108,c108,p12[6]);
	fa f147(s118,c119,s109,c109,p12[7]);
	fa f148(s119,c1110,s1010,c1010,p12[8]);
	fa f149(s1110,c1111,s1011,c1011,p12[9]);
	fa f150(s1111,c1112,s1012,c1012,p12[10]);
	fa f151(s1112,c1113,s1013,c1013,p12[11]);
	fa f152(s1113,c1114,s1014,c1014,p12[12]);
	fa f153(s1114,c1115,s1015,c1015,p12[13]);
	fa h22(s1115,c1116,p11[15],p12[14],c1016);
	//stage12
	ha h23(out1[12],c121,s11_1,c11_1);
	fa f154(s121,c122,s11_2,c11_2,p13[0]);
	fa f155(s122,c123,s11_3,c11_3,p13[1]);
	fa f156(s123,c124,s11_4,c11_4,p13[2]);
	fa f157(s124,c125,s11_5,c11_5,p13[3]);
	fa f158(s125,c126,s116,c11_6,p13[4]);
	fa f159(s126,c127,s117,c117,p13[5]);
	fa f160(s127,c128,s118,c118,p13[6]);
	fa f161(s128,c129,s119,c119,p13[7]);
	fa f162(s129,c1210,s1110,c1110,p13[8]);
	fa f163(s1210,c1211,s1111,c1111,p13[9]);
	fa f164(s1211,c1212,s1112,c1112,p13[10]);
	fa f165(s1212,c1213,s1113,c1113,p13[11]);
	fa f166(s1213,c1214,s1114,c1114,p13[12]);
	fa f167(s1214,c1215,s1115,c1115,p13[13]);
	fa h24(s1215,c1216,p12[15],p13[14],c1116);
	//stage13
	ha h25(out1[13],c131,s121,c121);
	fa f168(s131,c132,s122,c122,p14[0]);
	fa f169(s132,c133,s123,c123,p14[1]);
	fa f170(s133,c134,s124,c124,p14[2]);
	fa f171(s134,c135,s125,c125,p14[3]);
	fa f172(s135,c136,s126,c126,p14[4]);
	fa f173(s136,c137,s127,c127,p14[5]);
	fa f1700(s137,c138,s128,c128,p14[6]);
	fa f1741(s138,c139,s129,c129,p14[7]);
	fa f175(s139,c1310,s1210,c1210,p14[8]);
	fa f176(s1310,c1311,s1211,c1211,p14[9]);
	fa f177(s1311,c1312,s1212,c1212,p14[10]);
	fa f178(s1312,c1313,s1213,c1213,p14[11]);
	fa f179(s1313,c1314,s1214,c1214,p14[12]);
	fa f180(s1314,c1315,s1215,c1215,p14[13]);
	fa h26(s1315,c1316,p13[15],p14[14],c1216);
	
	//stage14
	ha h27(out1[14],c141,s131,c131);
	fa f181(s141,c142,s132,c132,p15[0]);
	fa f182(s142,c143,s133,c133,p15[1]);
	fa f183(s143,c144,s134,c134,p15[2]);
	fa f184(s144,c145,s135,c135,p15[3]);
	fa f185(s145,c146,s136,c136,p15[4]);
	fa f186(s146,c147,s137,c137,p15[5]);
	fa f187(s147,c148,s138,c138,p15[6]);
	fa f1881(s148,c149,s139,c139,p15[7]);
	fa f189(s149,c1410,s1310,c1310,p15[8]);
	fa f190(s1410,c1411,s1311,c1311,p15[9]);
	fa f191(s1411,c1412,s1312,c1312,p15[10]);
	fa f192(s1412,c1413,s1313,c1313,p15[11]);
	fa f193(s1413,c1414,s1314,c1314,p15[12]);
	fa f194(s1414,c1415,s1315,c1315,p15[13]);
	fa h28(s1415,c1416,p14[15],p15[14],c1316);
	
	//stage15
	ha h88(out1[15],cc1,s141,c141);
	fa h29(out2[0],c151,s142,c142,cc1);
	fa h30(out2[1],c152,s143,c143,c151);
	fa h31(out2[2],c153,s144,c144,c152);
	fa h32(out2[3],c154,s145,c145,c153);
	fa h33(out2[4],c155,s146,c146,c154);
	fa h34(out2[5],c156,s147,c147,c155);
	fa h35(out2[6],c157,s148,c148,c156);
	fa h36(out2[7],c158,s149,c149,c157);
	fa h37(out2[8],c159,s1410,c1410,c158);
	fa h38(out2[9],c1510,s1411,c1411,c159);
	fa h39(out2[10],c1511,s1412,c1412,c1510);
	fa h40(out2[11],c1512,s1413,c1413,c1511);
	fa h41(out2[12],c1513,s1414,c1414,c1512);
	fa h42(out2[13],c1514,s1415,c1415,c1513);
	fa hk(out2[14],c1515,s1415,c1416,c1514);
	ha h45(out2[15],c1516,p15[15],c1515);
	
	
	assign of=c1516;
	 
	 
	 

	 
endmodule
module fa(s,cout,A,cin,B);
input A,B,cin;
output s,cout;
wire s1,c1,c2;
xor g1(s1,A,B),g2(s,s1,cin),
	g3(cout,c2,c1);
	and g4(c1,A,B),g5(c2,s1,cin);
endmodule

module ha(S,Cout,in1,in2);
input in1,in2;
output S,Cout;
xor g6(S,in1,in2);
and g7(Cout,in1,in2);
endmodule
